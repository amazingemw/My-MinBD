module pipeline_two_tb();

reg [10:0] nty;  
reg [10:0] sty; 
reg [10:0] ety; 
reg [10:0] wty;
reg clk;
wire [10:0] nxt;
wire [10:0] sxt;
wire [10:0] ext;
wire [10:0] wxt;

always begin
#5.5 clk = ~clk;
end

initial begin
    clk = 0;	
    nty = 11'bz;
    sty = 11'b0000000101;
    ety = 11'b1000100001;
    wty = 11'b0000100100;

#5 nty = 11'b1000100100; //l
    sty = 11'b0000111111; //e
    ety = 11'b0000101100; //n
    wty = 11'b0000011100; //w

#5 nty = 11'b0000100110; //e
    sty = 11'b0000000001; //w
    ety = 11'b1000101100; //l
    wty = 11'b0000100100; //w

#5  nty = 11'b0000111100; //n
    sty = 11'b0000000011; //w
    ety = 11'b0000100100; //s
    wty = 11'b0000010101; //e

#5 nty = 11'b0000100100; //w
    sty = 11'b0000110100; //n
    ety = 11'bz; //e
    wty = 11'b0000100111; //l

end


pipeline_two U0 (
nty,
sty,
ety,
wty,
clk,
nxt,
sxt,
ext,
wxt
);


endmodule
